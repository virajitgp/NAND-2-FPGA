module RAM16K(
    input wire clk,             // Clock input
    input wire load,            // Write enable
    input wire [13:0] address,  // 14-bit address (0-16383)
    input wire [15:0] in,       // 16-bit input data
    output reg [15:0] out       // 16-bit output data
);
    // 16384 registers, each 16-bit wide
    reg [15:0] memory [0:16383];
    


    // Write operation
    always @(posedge clk) begin
        if (load) begin
            memory[address] <= in;
        end
    end

    // Read operation (update on address change)
    always @(posedge) begin
        out = memory[address];
    end

endmodule

